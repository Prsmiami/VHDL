library ieee;use ieee.std_logic_1164.all;Entity TriStateBuffer8 is  Port(Data : in std_logic_vector(7 downto 0);       En : in std_logic;       Outp1 : out std_logic_vector(15 downto 0));end;Architecture behav of TriStateBuffer8 is  begin    process(Data, En)      begin      if (En = '1') then        Outp1(7 downto 0) <= Data;
				Outp1(15 downto 8) <= "00000000";      else        Outp1 <= "ZZZZZZZZZZZZZZZZ";      end if;    end process;end behav;
