
module pll (
	clk_clk,
	reset_1_reset_n,
	clk_in_clk,
	clk_out_clk,
	reset_reset);	

	input		clk_clk;
	input		reset_1_reset_n;
	input		clk_in_clk;
	output		clk_out_clk;
	input		reset_reset;
endmodule
