library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity loop_counter is
  
port( cntr_in: IN std_logic_vector(13 downto 0); --Data input
      clk,load: IN std_logic; --Clock
			CE: OUT std_logic ; --Counter Expired signal
      cntr_out: OUT std_logic_vector(13 downto 0) --Data output     
 );
end loop_counter;

architecture behav of loop_counter is
	signal count : integer;
	signal Reg1 : integer;   	 
begin
  process(clk) -- Do this every time the clock changes
  begin
      CE <= '0';
    if (load = '1') then
     	count<=conv_integer(cntr_in);
	elsif (count <= 1) then
     	CE<='1';
    elsIf (clk = '1' and clk' event) then
		Reg1 <= count-1;
   		count <= Reg1;
    end if ;
    cntr_out <= cntr_in; --conv_std_logic_vector(count, 14); 
	end process;
end behav;
